`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    05:03:51 10/05/2021 
// Design Name: 
// Module Name:    MSDAP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module main(
    output reg [39:0] dataOut,
    input clk,
    input rst
    );
    
    reg [15:0] coeff = {
        16'h00BF,      // 1
        16'h015A,      // 2
        16'h01CE,      // 3
        16'h014C,      // 4
        16'h00D5,      // 5
        16'h015E,      // 6
        16'h01F1,      // 7
        16'h011D,      // 8
        16'h0051,      // 9
        16'h0141,      // 10
        16'h014D,      // 11
        16'h0056,      // 12
        16'h0092,      // 13
        16'h01E0,      // 14
        16'h0161,      // 15
        16'h011A,      // 16
        16'h0018,      // 17
        16'h016E,      // 18
        16'h01B3,      // 19
        16'h005F,      // 20
        16'h00DD,      // 21
        16'h0071,      // 22
        16'h0157,      // 23
        16'h0024,      // 24
        16'h01F7,      // 25
        16'h00C9,      // 26
        16'h00D0,      // 27
        16'h0054,      // 28
        16'h01CC,      // 29
        16'h00D8,      // 30
        16'h004B,      // 31
        16'h00D3,      // 32
        16'h018A,      // 33
        16'h00E0,      // 34
        16'h017D,      // 35
        16'h01E4,      // 36
        16'h010F,      // 37
        16'h008D,      // 38
        16'h004F,      // 39
        16'h0160,      // 40
        16'h0101,      // 41
        16'h0047,      // 42
        16'h0158,      // 43
        16'h0183,      // 44
        16'h010B,      // 45
        16'h01FA,      // 46
        16'h00E5,      // 47
        16'h0184,      // 48
        16'h01FB,      // 49
        16'h0124,      // 50
        16'h012B,      // 51
        16'h00B2,      // 52
        16'h013A,      // 53
        16'h00B3,      // 54
        16'h0011,      // 55
        16'h0012,      // 56
        16'h0171,      // 57
        16'h0157,      // 58
        16'h003E,      // 59
        16'h0043,      // 60
        16'h0026,      // 61
        16'h00BC,      // 62
        16'h0175,      // 63
        16'h00F8,      // 64
        16'h00EB,      // 65
        16'h001A,      // 66
        16'h00BD,      // 67
        16'h0017,      // 68
        16'h00D2,      // 69
        16'h01A7,      // 70
        16'h00A6,      // 71
        16'h007F,      // 72
        16'h0161,      // 73
        16'h01A3,      // 74
        16'h0064,      // 75
        16'h0118,      // 76
        16'h0076,      // 77
        16'h00CA,      // 78
        16'h00D0,      // 79
        16'h01B6,      // 80
        16'h0149,      // 81
        16'h01D7,      // 82
        16'h014C,      // 83
        16'h01C3,      // 84
        16'h00ED,      // 85
        16'h0194,      // 86
        16'h012F,      // 87
        16'h00E3,      // 88
        16'h0074,      // 89
        16'h01BD,      // 90
        16'h01C7,      // 91
        16'h0143,      // 92
        16'h0121,      // 93
        16'h003C,      // 94
        16'h017B,      // 95
        16'h0109,      // 96
        16'h0014,      // 97
        16'h0138,      // 98
        16'h00FE,      // 99
        16'h01F2,      // 100
        16'h0049,      // 101
        16'h011A,      // 102
        16'h01A4,      // 103
        16'h011D,      // 104
        16'h0059,      // 105
        16'h006A,      // 106
        16'h015D,      // 107
        16'h01C8,      // 108
        16'h007E,      // 109
        16'h01FA,      // 110
        16'h00A0,      // 111
        16'h01BE,      // 112
        16'h0083,      // 113
        16'h01E2,      // 114
        16'h018B,      // 115
        16'h00E2,      // 116
        16'h01C8,      // 117
        16'h005F,      // 118
        16'h0003,      // 119
        16'h0172,      // 120
        16'h0013,      // 121
        16'h0073,      // 122
        16'h01C4,      // 123
        16'h01D2,      // 124
        16'h01A4,      // 125
        16'h001F,      // 126
        16'h013D,      // 127
        16'h0030,      // 128
        16'h009E,      // 129
        16'h017A,      // 130
        16'h0199,      // 131
        16'h0011,      // 132
        16'h01CD,      // 133
        16'h0083,      // 134
        16'h0128,      // 135
        16'h0076,      // 136
        16'h01E1,      // 137
        16'h0029,      // 138
        16'h01FF,      // 139
        16'h0160,      // 140
        16'h00B5,      // 141
        16'h0180,      // 142
        16'h0077,      // 143
        16'h0150,      // 144
        16'h0051,      // 145
        16'h01CC,      // 146
        16'h00AC,      // 147
        16'h0030,      // 148
        16'h01DE,      // 149
        16'h004A,      // 150
        16'h01AC,      // 151
        16'h00E2,      // 152
        16'h01D3,      // 153
        16'h0052,      // 154
        16'h001E,      // 155
        16'h01C6,      // 156
        16'h01ED,      // 157
        16'h00CD,      // 158
        16'h01AA,      // 159
        16'h0065,      // 160
        16'h0199,      // 161
        16'h0012,      // 162
        16'h00E7,      // 163
        16'h00D6,      // 164
        16'h0148,      // 165
        16'h0192,      // 166
        16'h00E8,      // 167
        16'h0015,      // 168
        16'h0176,      // 169
        16'h01B6,      // 170
        16'h0026,      // 171
        16'h01CC,      // 172
        16'h01DA,      // 173
        16'h004C,      // 174
        16'h0067,      // 175
        16'h0174,      // 176
        16'h000C,      // 177
        16'h01D7,      // 178
        16'h00D8,      // 179
        16'h01E9,      // 180
        16'h010A,      // 181
        16'h01DE,      // 182
        16'h0157,      // 183
        16'h01D4,      // 184
        16'h00AE,      // 185
        16'h00FB,      // 186
        16'h0110,      // 187
        16'h00E4,      // 188
        16'h0099,      // 189
        16'h0019,      // 190
        16'h01C2,      // 191
        16'h0122,      // 192
        16'h0163,      // 193
        16'h0006,      // 194
        16'h0068,      // 195
        16'h01C6,      // 196
        16'h01D0,      // 197
        16'h00DB,      // 198
        16'h011B,      // 199
        16'h0152,      // 200
        16'h01D1,      // 201
        16'h0084,      // 202
        16'h017A,      // 203
        16'h0111,      // 204
        16'h0096,      // 205
        16'h0046,      // 206
        16'h01CA,      // 207
        16'h009C,      // 208
        16'h0168,      // 209
        16'h010F,      // 210
        16'h0110,      // 211
        16'h00C7,      // 212
        16'h00C8,      // 213
        16'h0181,      // 214
        16'h0149,      // 215
        16'h0124,      // 216
        16'h017D,      // 217
        16'h01F0,      // 218
        16'h01F3,      // 219
        16'h0030,      // 220
        16'h014D,      // 221
        16'h01BA,      // 222
        16'h01D2,      // 223
        16'h01B2,      // 224
        16'h0161,      // 225
        16'h01BC,      // 226
        16'h0120,      // 227
        16'h01DD,      // 228
        16'h01B3,      // 229
        16'h0166,      // 230
        16'h01D7,      // 231
        16'h00CB,      // 232
        16'h00D5,      // 233
        16'h01A2,      // 234
        16'h0107,      // 235
        16'h0173,      // 236
        16'h0032,      // 237
        16'h017B,      // 238
        16'h0151,      // 239
        16'h00E9,      // 240
        16'h0123,      // 241
        16'h0082,      // 242
        16'h0075,      // 243
        16'h0057,      // 244
        16'h015B,      // 245
        16'h001A,      // 246
        16'h00C3,      // 247
        16'h013E,      // 248
        16'h01D8,      // 249
        16'h00A7,      // 250
        16'h00C4,      // 251
        16'h00D3,      // 252
        16'h00E7,      // 253
        16'h00CD,      // 254
        16'h018E,      // 255
        16'h01A1,      // 256
        16'h012E,      // 257
        16'h00D2,      // 258
        16'h0116,      // 259
        16'h013D,      // 260
        16'h01FA,      // 261
        16'h0180,      // 262
        16'h017A,      // 263
        16'h005F,      // 264
        16'h002E,      // 265
        16'h015A,      // 266
        16'h00F9,      // 267
        16'h0067,      // 268
        16'h0150,      // 269
        16'h012C,      // 270
        16'h00AD,      // 271
        16'h01D4,      // 272
        16'h0089,      // 273
        16'h000D,      // 274
        16'h011C,      // 275
        16'h01EF,      // 276
        16'h007B,      // 277
        16'h00DC,      // 278
        16'h015E,      // 279
        16'h01A8,      // 280
        16'h015B,      // 281
        16'h005C,      // 282
        16'h0038,      // 283
        16'h01CC,      // 284
        16'h0137,      // 285
        16'h019E,      // 286
        16'h00E5,      // 287
        16'h00B2,      // 288
        16'h01C7,      // 289
        16'h016E,      // 290
        16'h0003,      // 291
        16'h018C,      // 292
        16'h00B7,      // 293
        16'h009C,      // 294
        16'h00C1,      // 295
        16'h0045,      // 296
        16'h019E,      // 297
        16'h0022,      // 298
        16'h0029,      // 299
        16'h0167,      // 300
        16'h00C5,      // 301
        16'h0177,      // 302
        16'h014F,      // 303
        16'h0033,      // 304
        16'h012E,      // 305
        16'h012B,      // 306
        16'h01BB,      // 307
        16'h01C9,      // 308
        16'h00AF,      // 309
        16'h010F,      // 310
        16'h00BD,      // 311
        16'h0113,      // 312
        16'h01B8,      // 313
        16'h01F0,      // 314
        16'h0150,      // 315
        16'h01DF,      // 316
        16'h008F,      // 317
        16'h0030,      // 318
        16'h0177,      // 319
        16'h01D3,      // 320
        16'h0009,      // 321
        16'h017F,      // 322
        16'h0072,      // 323
        16'h0031,      // 324
        16'h007A,      // 325
        16'h016D,      // 326
        16'h010B,      // 327
        16'h013C,      // 328
        16'h0065,      // 329
        16'h01CC,      // 330
        16'h0123,      // 331
        16'h01AD,      // 332
        16'h01F6,      // 333
        16'h0044,      // 334
        16'h0073,      // 335
        16'h01AB,      // 336
        16'h0029,      // 337
        16'h01D4,      // 338
        16'h01EF,      // 339
        16'h0080,      // 340
        16'h00E0,      // 341
        16'h00F0,      // 342
        16'h01C8,      // 343
        16'h01B3,      // 344
        16'h009B,      // 345
        16'h00F2,      // 346
        16'h0142,      // 347
        16'h00C5,      // 348
        16'h018A,      // 349
        16'h00A6,      // 350
        16'h01B5,      // 351
        16'h0147,      // 352
        16'h0094,      // 353
        16'h00AE,      // 354
        16'h0051,      // 355
        16'h018B,      // 356
        16'h018C,      // 357
        16'h019C,      // 358
        16'h008D,      // 359
        16'h01E8,      // 360
        16'h00FB,      // 361
        16'h0112,      // 362
        16'h0033,      // 363
        16'h011E,      // 364
        16'h01B6,      // 365
        16'h01DD,      // 366
        16'h00B1,      // 367
        16'h019C,      // 368
        16'h0071,      // 369
        16'h0124,      // 370
        16'h00DB,      // 371
        16'h01E4,      // 372
        16'h00A9,      // 373
        16'h00ED,      // 374
        16'h01B9,      // 375
        16'h0020,      // 376
        16'h002F,      // 377
        16'h0199,      // 378
        16'h0075,      // 379
        16'h0034,      // 380
        16'h009D,      // 381
        16'h00A8,      // 382
        16'h0068,      // 383
        16'h0014,      // 384
        16'h01BE,      // 385
        16'h00D4,      // 386
        16'h01D6,      // 387
        16'h017B,      // 388
        16'h0017,      // 389
        16'h01B2,      // 390
        16'h014C,      // 391
        16'h0143,      // 392
        16'h0126,      // 393
        16'h00E1,      // 394
        16'h0191,      // 395
        16'h01F9,      // 396
        16'h00A0,      // 397
        16'h01D1,      // 398
        16'h01CA,      // 399
        16'h00D5,      // 400
        16'h0051,      // 401
        16'h0007,      // 402
        16'h00BF,      // 403
        16'h015A,      // 404
        16'h01CE,      // 405
        16'h014C,      // 406
        16'h00D5,      // 407
        16'h015E,      // 408
        16'h01F1,      // 409
        16'h011D,      // 410
        16'h0051,      // 411
        16'h0141,      // 412
        16'h014D,      // 413
        16'h0056,      // 414
        16'h0092,      // 415
        16'h01E0,      // 416
        16'h0161,      // 417
        16'h011A,      // 418
        16'h0018,      // 419
        16'h016E,      // 420
        16'h01B3,      // 421
        16'h005F,      // 422
        16'h00DD,      // 423
        16'h0071,      // 424
        16'h0157,      // 425
        16'h0024,      // 426
        16'h01F7,      // 427
        16'h00C9,      // 428
        16'h00D0,      // 429
        16'h0054,      // 430
        16'h01CC,      // 431
        16'h00D8,      // 432
        16'h004B,      // 433
        16'h00D3,      // 434
        16'h018A,      // 435
        16'h00E0,      // 436
        16'h017D,      // 437
        16'h01E4,      // 438
        16'h010F,      // 439
        16'h008D,      // 440
        16'h004F,      // 441
        16'h0160,      // 442
        16'h0101,      // 443
        16'h0047,      // 444
        16'h0158,      // 445
        16'h0183,      // 446
        16'h010B,      // 447
        16'h01FA,      // 448
        16'h00E5,      // 449
        16'h0184,      // 450
        16'h01FB,      // 451
        16'h0124,      // 452
        16'h012B,      // 453
        16'h00B2,      // 454
        16'h013A,      // 455
        16'h00B3,      // 456
        16'h0011,      // 457
        16'h0012,      // 458
        16'h0171,      // 459
        16'h0157,      // 460
        16'h003E,      // 461
        16'h0043,      // 462
        16'h0026,      // 463
        16'h00BC,      // 464
        16'h0175,      // 465
        16'h00F8,      // 466
        16'h00EB,      // 467
        16'h001A,      // 468
        16'h00BD,      // 469
        16'h0017,      // 470
        16'h00D2,      // 471
        16'h01A7,      // 472
        16'h00A6,      // 473
        16'h007F,      // 474
        16'h0161,      // 475
        16'h01A3,      // 476
        16'h0064,      // 477
        16'h0118,      // 478
        16'h0076,      // 479
        16'h00CA,      // 480
        16'h00D0,      // 481
        16'h01B6,      // 482
        16'h0149,      // 483
        16'h01D7,      // 484
        16'h014C,      // 485
        16'h01C3,      // 486
        16'h00ED,      // 487
        16'h0194,      // 488
        16'h012F,      // 489
        16'h00E3,      // 490
        16'h0074,      // 491
        16'h01BD,      // 492
        16'h01C7,      // 493
        16'h0143,      // 494
        16'h0121,      // 495
        16'h003C,      // 496
        16'h017B,      // 497
        16'h0109,      // 498
        16'h0014,      // 499
        16'h0138,      // 500
        16'h00FE,      // 501
        16'h01F2,      // 502
        16'h0049,      // 503
        16'h011A,      // 504
        16'h01A4,      // 505
        16'h011D,      // 506
        16'h0059,      // 507
        16'h006A,      // 508
        16'h015D,      // 509
        16'h01C8,      // 510
        16'h007E,      // 511
        16'h01FA       // 512
    };
    
    reg [7:0] rj = {
        8'h0020,      // r1
        8'h0020,      // r2
        8'h0020,      // r3
        8'h0020,      // r4
        8'h0020,      // r5
        8'h0020,      // r6
        8'h0020,      // r7
        8'h0020,      // r8
        8'h0020,      // r9
        8'h0020,      // r10
        8'h0020,      // r11
        8'h0020,      // r12
        8'h0020,      // r13
        8'h0020,      // r14
        8'h0020,      // r15
        8'h0020      // r16
    };
    
//    reg [15:0] data = {
//        16'hC48B,
//        16'hCEAD,
//        16'hC747,
//        16'h93B7,
//        16'hDDA7,
//        16'hC760,
//        16'h5DFC,
//        16'h8817,
//        16'h86D8,
//        16'h3498,
//        16'hB570,
//        16'h366E,
//        16'hDB45,
//        16'h20B6,
//        16'h2F04,
//        16'hFB27,
//        16'h20AA,
//        16'hDA4F,
//        16'h8EEB,
//        16'hB61F,
//        16'h39D5,
//        16'h75AA,
//        16'h7AB1,
//        16'h4C2A,
//        16'h312A,
//        16'h4744,
//        16'hFEB1,
//        16'h268D,
//        16'hB41F,
//        16'h6B4C,
//        16'h0A9C,
//        16'hB182,
//        16'h94C0,
//        16'h3F27,
//        16'hF2F9,
//        16'hDDB7,
//        16'h482D,
//        16'hE7ED,
//        16'hEEA0,
//        16'h9FCE,
//        16'h6817,
//        16'hC7EA,
//        16'h983E,
//        16'h70DF,
//        16'h3247,
//        16'h0D1E,
//        16'h71D4,
//        16'hCBF2,
//        16'h0817,
//        16'h25BE,
//        16'h5C37,
//        16'hB286,
//        16'hF0F6,
//        16'h42B0,
//        16'h2092,
//        16'h2A0C,
//        16'h13E8,
//        16'hDC13,
//        16'hEBDF,
//        16'hBB6C,
//        16'h3E04,
//        16'h2DB5,
//        16'hCA72,
//        16'hF17F
//    };

    //Integers, equivalent to signed 32 bit register: reg signed [31:0]
    integer n, j, i, prevRj, dataIndex, endPoint;
    integer dataSize; // = 64;
    integer rjSize = 16;
    
    //Registers
    reg [39:0] overallResult, currentResult;
    reg coeffSign, sign;
    reg [8:0] tempCoeff;
    reg [7:0] coeffValue;
    reg [23:0] dataX;
    reg [23:0] tempDataX;
    reg [39:0] ujTemp = 0; 
    reg [39:0] tempData;
    
    //Instantiate memory module
    rom memory(.clk(clk), .address(dataIndex), .data(dataX));
    
    always @ (posedge clk) begin
    
        // Main loop. needs dataSize from input file
        for(n = 0; n < dataSize; n = n + 1) begin
            overallResult = 0;
            prevRj = 0;
        
            // Second loop in main function
            for(j = 0; j < rjSize; j = j + 1) begin
            
                currentResult = 0;
                endPoint = prevRj + rj[j];  //Pre-calculate value of prevRj + rj[j]
                
                // Calculate Uj Fucntion ---------------------------------------------------------------------------------------------------------------
                for (i = prevRj; i < endPoint; i = i + 1) begin
                    
                    tempCoeff = coeff[i];           //Get currrent coefficient from memory array
                    coeffSign = tempCoeff[1];       //Extract sign
                    coeffValue = tempCoeff[7:0];    //Extract value
                    
                    dataIndex = n - coeffValue;     //Calculate index of data to retrieve, this is an input to the rom module,
                                                    //and will tell the rom what address to retrieve data from
                    if(dataIndex < 0) begin         // If index is lesss than zero, result is 0
                        ujTemp = ujTemp + 0;
                    end
                    else begin

                        //dataX = data[dataIndex];
                        sign = dataX[15];           //dataX is the output from rom, represents the data retrieved from rom.
                                                    //Note that output from rom is 16 bits, and dataX is 24 bits.

                        if(sign) begin
			                 tempDataX = dataX | 'hFF0000;   //Pad with 1's if negative
		                end
		                else begin
			                 tempDataX = dataX & 'h00FFFF;   //Pad with 0's if positive
		                end
                        
                        if(coeffSign == 1) begin
                            tempData = {((~tempDataX) + 1), 16'h000};   //Twos compliment if negative. Then set the most significant 24 bits to contain data
                                                                        //tempData is 40 bits, tempDataX is 24 bits. The most significant 24bits are occupied
                                                                        //by tempDataX and the 16 LSBs are filled with 0's
                            ujTemp = ujTemp + tempData;                 //Add to running total
                        end
                        else begin
                            tempData = {tempDataX, 16'h0000};           //If positive, just set most significant bits to hold data.
                            ujTemp = ujTemp + tempData;                 //Add to running total
                        end
                    end
                    
                end
            
                currentResult = ujTemp;                                 //Set current result to final total
                // --------------------------------------------------------------------------------------------------------------------------------
                
                overallResult = overallResult + currentResult;          //Add to running total
                
                //This is equivalwent to the shiftResultRight1Bit function.
                if(overallResult[39] == 1) begin
                    overallResult = (overallResult >> 1) | 'h8000000000; //If negative, shift right and pad with 1
                end
                else begin
                    overallResult = overallResult >> 1;                 //If positive, shift right and pad with 0
                end
                
                prevRj = endPoint;      //endpoint was set to prevRj + rj[j] at the beginning of the loop.
            
            end
            
            dataOut = overallResult; // >> 24; not sure if we need this shift operation here.
        
        end
    
    end

endmodule
