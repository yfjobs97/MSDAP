`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    05:14:41 10/05/2021 
// Design Name: 
// Module Name:    calculateUj 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module calculateUj(
    input n,
    input [23:0] dataX,
    input [8:0] coeff,
    input startPoint,
    input endPoint,
    output uj
    );


endmodule
