`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    05:03:51 10/05/2021 
// Design Name: 
// Module Name:    MSDAP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module main(
    output [39:0] dataOut,
    input [15:0] dataIn,
    input [11:0] coeff,
    input [8:0] rj
    );


endmodule
